LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Testbench_Adder4BitParity IS
END ENTITY;

ARCHITECTURE Testbench OF Testbench_Adder4BitParity IS


	-- Signale fuer die Eingabe- und Ausgabewerte
	SIGNAL A, B : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL SUM : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL EVEN_PARITY, ODD_PARITY : BIT;
    
    -- Signals Testbench
	SIGNAL SUM_XNOR_DESIRED_CONDITION4, 
           SUM_XNOR_DESIRED_CONDITION3, 
           SUM_XNOR_DESIRED_CONDITION2, 
           SUM_XNOR_DESIRED_CONDITION1, 
           SUM_XNOR_DESIRED_CONDITION0 : STD_LOGIC;
    SIGNAL EVEN_PARITY_DESIRED_CONDITION, 
           ODD_PARITY_DESIRED_CONDITION, 
           EVEN_PARITY_XNOR_DESIRED_CONDITION, 
           ODD_PARITY_XNOR_DESIRED_CONDITION : BIT;
	SIGNAL SUM_DESIRED_CONDITION : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN
	DUT: ENTITY WORK.Adder4BitParity
		PORT MAP (
			A => A,
			B => B,
			SUM => SUM,
			EVEN_PARITY => EVEN_PARITY,
			ODD_PARITY => ODD_PARITY
		);

	-- Testprozess
	PROCESS
	BEGIN
		-- Testfall 1: Hoechster Zustand
		SUM_DESIRED_CONDITION <= "11110";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "1111";
		B <= "1111";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
        
		-- Testfall 2: Kleinster Zustand
		SUM_DESIRED_CONDITION <= "00000";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "0000";
		B <= "0000";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
        
		-- Testfall 3: Zustand dazwischen 1
		SUM_DESIRED_CONDITION <= "00001";
        EVEN_PARITY_DESIRED_CONDITION <= '1';
        ODD_PARITY_DESIRED_CONDITION <= '0';
		
		A <= "0001";
		B <= "0000";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
        
		-- Testfall 4: Zustand dazwischen 2
		SUM_DESIRED_CONDITION <= "01111";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "1001";
		B <= "0110";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
		
		-- Testfall 5: Zustand dazwischen 3
		SUM_DESIRED_CONDITION <= "11011";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "1101";
		B <= "1110";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
        
		-- Testfall 6: Zustand dazwischen 4
		SUM_DESIRED_CONDITION <= "10101";
        EVEN_PARITY_DESIRED_CONDITION <= '1';
        ODD_PARITY_DESIRED_CONDITION <= '0';
		
		A <= "1110";
		B <= "0111";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;

		-- Testfall 7: Zustand dazwischen 5
		SUM_DESIRED_CONDITION <= "10001";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "0101";
		B <= "1100";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
		
		-- Testfall 8: Zustand dazwischen 6
		SUM_DESIRED_CONDITION <= "00101";
        EVEN_PARITY_DESIRED_CONDITION <= '0';
        ODD_PARITY_DESIRED_CONDITION <= '1';
		
		A <= "0001";
		B <= "0100";
		WAIT FOR 0.1 ns;
		SUM_XNOR_DESIRED_CONDITION4 <= SUM(4) XNOR SUM_DESIRED_CONDITION(4); -- I
        SUM_XNOR_DESIRED_CONDITION3 <= SUM(3) XNOR SUM_DESIRED_CONDITION(3); -- HATE
        SUM_XNOR_DESIRED_CONDITION2 <= SUM(2) XNOR SUM_DESIRED_CONDITION(2); -- YOU
        SUM_XNOR_DESIRED_CONDITION1 <= SUM(1) XNOR SUM_DESIRED_CONDITION(1);
        SUM_XNOR_DESIRED_CONDITION0 <= SUM(0) XNOR SUM_DESIRED_CONDITION(0);
        
        EVEN_PARITY_XNOR_DESIRED_CONDITION <= EVEN_PARITY XNOR EVEN_PARITY_DESIRED_CONDITION;
        ODD_PARITY_XNOR_DESIRED_CONDITION <= ODD_PARITY XNOR ODD_PARITY_DESIRED_CONDITION;
		WAIT FOR 10 ns;
		
		-- Hier koennen weitere Testfaelle hinzugefuegt werden
        
		WAIT; -- Endlosschleife
	END PROCESS;
END ARCHITECTURE;

